/*
    This sprite table was generated using 'conv_to_sv.py'. Find out more here: https://github.com/Atrifex/ECE385-HelperTools
    To use, instantiate this module in your color mapper. The SpriteX input should be connected to
        'ObjectXSize - DistX', where ObjectXSize is the width of your object in pixels along the
        x direction. DistX is the horizontal distance between the DrawX pxiel and the top left corner
        of the object in question, so something like: 'DistX = DrawX - ObjectXPosition' is fine.
        Similarly this goes for SpriteY. Warning: If you don't do this, your image will be flipped along
        the axis you ignored. This is a handy way to flip an image if you need to, though.
 
    In the color mapper, you can then simply do something like:
    module ColorMapper(...)
    ...
    logic [7:0] ObjectR, ObjectG, ObjectB
    parameter ObjectXSize = 10'd10;
    ...
    always_comb
    ...
         if(ObjectOn == 1'b1)
         begin
             Red = ObjectR
             Green = ObjectG
             Blue = ObjectB
         end
     ...
     ObjectSpriteTable ost(
                           .SpriteX(ObjectXSize - DistX), .SpriteY(ObjectYSize - DistY),
                           .SpriteR(ObjectR), .SpriteG(ObjectG), .SpriteB(ObjectB)
                           );
 
     See the comment at the top of the generation script if you're still confused.
*/
module GameOver(input [9:0] SpriteX, SpriteY,
            output [7:0] SpriteR, SpriteG, SpriteB);

parameter bit [7:0] SpritePaletteR[6:0] = '{8'd0, 8'd144, 8'd182, 8'd102, 8'd58, 8'd219, 8'd255};

parameter bit [2:0] SpriteTableR[14:0][140:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd4,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0},
'{3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0},
'{3'd0,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd5,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd2,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd6,3'd6,3'd6,3'd4,3'd0,3'd3,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0},
'{3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd0,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd5,3'd6,3'd6,3'd1,3'd0,3'd2,3'd6,3'd6,3'd1,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0},
'{3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd2,3'd0,3'd2,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd1,3'd6,3'd6,3'd2,3'd0,3'd6,3'd6,3'd6,3'd4,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0},
'{3'd1,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd3,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd3,3'd6,3'd6,3'd6,3'd4,3'd6,3'd6,3'd6,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd1,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd6,3'd6,3'd6,3'd2,3'd6,3'd6,3'd2,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd5,3'd0,3'd5,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd4,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0},
'{3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd3,3'd4,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3}};

parameter bit [7:0] SpritePaletteG[6:0] = '{8'd0, 8'd144, 8'd102, 8'd182, 8'd58, 8'd219, 8'd255};

parameter bit [2:0] SpriteTableG[14:0][140:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0},
'{3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0},
'{3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd1,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd3,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd3,3'd6,3'd6,3'd5,3'd0,3'd0,3'd3,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0},
'{3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd3,3'd2,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd1,3'd6,3'd6,3'd6,3'd4,3'd0,3'd6,3'd6,3'd6,3'd1,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd5,3'd6,3'd6,3'd2,3'd2,3'd6,3'd6,3'd5,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd3,3'd6,3'd6,3'd3,3'd1,3'd6,3'd6,3'd3,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd5,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd2,3'd6,3'd6,3'd5,3'd5,3'd6,3'd6,3'd2,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd1,3'd4,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd5,3'd2,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0},
'{3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0},
'{3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd0,3'd1,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd5,3'd6,3'd6,3'd5,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0}};

parameter bit [7:0] SpritePaletteB[6:0] = '{8'd0, 8'd144, 8'd102, 8'd182, 8'd58, 8'd219, 8'd255};

parameter bit [2:0] SpriteTableB[14:0][140:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0},
'{3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0},
'{3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd3,3'd6,3'd6,3'd1,3'd0,3'd0,3'd6,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0},
'{3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd2,3'd3,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd1,3'd6,3'd6,3'd5,3'd0,3'd2,3'd6,3'd6,3'd5,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0},
'{3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd0,3'd2,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd4,3'd6,3'd6,3'd6,3'd0,3'd3,3'd6,3'd6,3'd1,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0},
'{3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd6,3'd6,3'd6,3'd2,3'd5,3'd6,3'd6,3'd2,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd5,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd3,3'd6,3'd6,3'd3,3'd6,3'd6,3'd6,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd1,3'd3,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd2,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd0,3'd1,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd5,3'd6,3'd6,3'd6,3'd0,3'd0,3'd4,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0,3'd0,3'd5,3'd6,3'd6,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd0}};

assign SpriteR = SpritePaletteR[SpriteTableR[SpriteY][SpriteX]];
assign SpriteG = SpritePaletteG[SpriteTableG[SpriteY][SpriteX]];
assign SpriteB = SpritePaletteB[SpriteTableB[SpriteY][SpriteX]];

endmodule
