module SpaceshipProjectileSprite(input [8:0] SpriteX, SpriteY,
            output [7:0] SpriteR, SpriteG, SpriteB);

