module GalagaText(input [9:0] SpriteX, SpriteY,
            output [7:0] SpriteR, SpriteG, SpriteB);

parameter bit [7:0] SpriteTableR[14:0][97:0] = '{'{8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hdb,8'h00,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hdb,8'h00,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00},
'{8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00},
'{8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00},
'{8'h90,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h66,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h66,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h66,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00},
'{8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00},
'{8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00},
'{8'h00,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00},
'{8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00},
'{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00},
'{8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66}};

parameter bit [7:0] SpriteTableG[14:0][97:0] = '{'{8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'h90,8'h00,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'h90,8'h00,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00},
'{8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hb6,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hb6,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hb6,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00},
'{8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00},
'{8'hdb,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00},
'{8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00},
'{8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00},
'{8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00},
'{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00},
'{8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00},
'{8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00}};

parameter bit [7:0] SpriteTableB[14:0][97:0] = '{'{8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'h3a,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'h3a,8'h3a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'h66,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'h66,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'h66,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'h00},
'{8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h00,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h00,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'h00,8'h66,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00},
'{8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00},
'{8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h00},
'{8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00},
'{8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'h66,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00},
'{8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00,8'h66,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h90,8'h00,8'h00},
'{8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdb,8'h00,8'h00},
'{8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hff,8'hff,8'hff,8'hff,8'h3a,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'hdb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h66,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00}};

assign SpriteR = SpriteTableR[SpriteY][SpriteX];
assign SpriteG = SpriteTableG[SpriteY][SpriteX];
assign SpriteB = SpriteTableB[SpriteY][SpriteX];

endmodule
