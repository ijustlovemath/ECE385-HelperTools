/*
    This sprite table was generated using 'conv_to_sv.py'. Find out more here: https://github.com/ijustlovemath/ECE385-HelperTools
    To use, instantiate this module in your color mapper. The SpriteX input should be connected to
        'ObjectXSize - DistX', where ObjectXSize is the width of your object in pixels along the
        x direction. DistX is the horizontal distance between the DrawX pxiel and the top left corner
        of the object in question, so something like: 'DistX = DrawX - ObjectXPosition' is fine.
        Similarly this goes for SpriteY. Warning: If you don't do this, your image will be flipped along
        the axis you ignored. This is a handy way to flip an image if you need to, though.
 
    In the color mapper, you can then simply do something like:
    module ColorMapper(...)
    ...
    logic [7:0] ObjectR, ObjectG, ObjectB
    parameter ObjectXSize = 10'd10;
    parameter ObjectYSize = 10'd10;
    ...
    always_comb
    ...
         if(ObjectOn == 1'b1)
         begin
             Red = ObjectR
             Green = ObjectG
             Blue = ObjectB
         end
     ...
     ObjectSpriteTable ost(
                           .SpriteX(ObjectXSize - DistX), .SpriteY(ObjectYSize - DistY),
                           .SpriteR(ObjectR), .SpriteG(ObjectG), .SpriteB(ObjectB)
                           );
 
     See the comment at the top of the generation script if you're still confused.
*/
module GalagaLogo(input [9:0] SpriteX, SpriteY,
            output [7:0] SpriteR, SpriteG, SpriteB);

logic [9:0] X_Index, Y_Index;

assign X_Index = SpriteX % 10'd32;
assign Y_Index = SpriteY % 10'd32;
logic [9:0] SpriteTableR;

parameter bit [7:0] SpritePaletteR[7:0] = '{8'd16, 8'd49, 8'd82, 8'd115, 8'd148, 8'd181, 8'd214, 8'd247};

	always_comb
	begin
		SpriteTableR = 10'd0;
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_31_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_31_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_31_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_31_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_30_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_30_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_30_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_30_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_29_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_29_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_29_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_29_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_28_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_28_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_28_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_28_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_27_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_27_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_27_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_27_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_26_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_26_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_26_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_26_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_25_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_25_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_25_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_25_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_24_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_24_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_24_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_24_28[Y_Index][X_Index];
		end
	end

parameter bit [2:0] SpriteTableR_31_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd4,3'd2,3'd3,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd6,3'd3,3'd2,3'd3,3'd4,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd7,3'd6,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd5,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd3,3'd6,3'd7}};

parameter bit [2:0] SpriteTableR_31_30[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd2,3'd3,3'd4,3'd4,3'd3,3'd2,3'd3,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd4,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd3,3'd6,3'd7,3'd7,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd4,3'd2,3'd3,3'd4,3'd4,3'd3,3'd2,3'd3,3'd6,3'd7,3'd7,3'd6,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd5,3'd2,3'd3,3'd4,3'd3,3'd4,3'd3,3'd2,3'd6,3'd7,3'd7,3'd6,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd5,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd6,3'd3,3'd3,3'd4,3'd3,3'd4,3'd3,3'd2,3'd4,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd7,3'd4,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd6,3'd7,3'd7,3'd5,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd7,3'd3,3'd3,3'd4,3'd3,3'd4,3'd4,3'd3,3'd2,3'd5,3'd7,3'd7,3'd6,3'd2,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd7,3'd7,3'd5,3'd2,3'd3,3'd4,3'd4,3'd3,3'd4,3'd3,3'd3,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd3,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd5,3'd2,3'd3,3'd4,3'd3,3'd4,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd2,3'd6,3'd7,3'd7,3'd3,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd6,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd5,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd6,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd6,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd5,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd6,3'd5,3'd5,3'd5,3'd5,3'd4,3'd5,3'd5},
'{3'd0,3'd1,3'd4,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd1,3'd1,3'd5,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd1,3'd1,3'd6,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd1,3'd6,3'd7,3'd7,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_31_29[31:0][31:0] = '{'{3'd1,3'd1,3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd6,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd5,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd2,3'd6,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5},
'{3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd6,3'd7},
'{3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd7,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd1,3'd1,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd1,3'd1,3'd1,3'd2,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_31_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_30_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd4,3'd2},
'{3'd1,3'd0,3'd1,3'd2,3'd4,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd4,3'd5,3'd6,3'd7,3'd6,3'd4,3'd3,3'd2,3'd3},
'{3'd1,3'd2,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd3,3'd3,3'd4,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd2,3'd3,3'd4,3'd3},
'{3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd5,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd7,3'd7,3'd5,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd5},
'{3'd5,3'd3,3'd2,3'd2,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd6,3'd7},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd2,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7},
'{3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd5},
'{3'd3,3'd3,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd7,3'd7,3'd7,3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1},
'{3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd3,3'd2,3'd5,3'd7,3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1},
'{3'd3,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd1,3'd1,3'd5,3'd7,3'd6,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd5,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd2,3'd1,3'd1,3'd1},
'{3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd3,3'd7,3'd7,3'd4,3'd3,3'd3,3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2}};

parameter bit [2:0] SpriteTableR_30_30[31:0][31:0] = '{'{3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd4,3'd7,3'd7,3'd3,3'd2,3'd2,3'd2,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd3},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd6,3'd7,3'd6,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd6,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd5,3'd6},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd5,3'd2,3'd5,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd3,3'd7,3'd7,3'd4,3'd5,3'd7,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd2,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd2,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd4,3'd7,3'd7,3'd7,3'd5,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd7,3'd7,3'd7,3'd6,3'd3,3'd4,3'd6,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd5,3'd7,3'd7,3'd6,3'd3,3'd2},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd6,3'd7,3'd7,3'd7,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd3,3'd2,3'd3,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd6,3'd7,3'd7,3'd5,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd3,3'd2,3'd4,3'd7,3'd7,3'd7,3'd5,3'd5,3'd6,3'd7},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd5,3'd7,3'd7,3'd5,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0,3'd2,3'd6,3'd7,3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd5,3'd7,3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd7,3'd4,3'd3,3'd3,3'd3,3'd4,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd7,3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd7,3'd7,3'd7,3'd3,3'd1,3'd0,3'd1,3'd5,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd5,3'd7,3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd5,3'd2,3'd0,3'd2,3'd7,3'd7},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd6,3'd7,3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd0,3'd3,3'd7,3'd7},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd6,3'd7,3'd7,3'd4,3'd1,3'd3,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd6,3'd2,3'd4,3'd7,3'd7},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd4,3'd5,3'd7,3'd6},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd6,3'd7,3'd7,3'd5},
'{3'd1,3'd0,3'd1,3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5},
'{3'd1,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd4},
'{3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd7,3'd7,3'd3},
'{3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd7,3'd7,3'd7,3'd2},
'{3'd6,3'd6,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd7,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd6,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd5,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd4,3'd0}};

parameter bit [2:0] SpriteTableR_30_29[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd7,3'd6,3'd1,3'd0},
'{3'd0,3'd1,3'd3,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd6,3'd6,3'd1,3'd0},
'{3'd2,3'd5,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd1,3'd1,3'd2,3'd6,3'd6,3'd1,3'd0},
'{3'd7,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd0,3'd1,3'd2,3'd6,3'd7,3'd3,3'd0},
'{3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd6,3'd3},
'{3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7},
'{3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd7},
'{3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd5},
'{3'd7,3'd6,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd7,3'd5,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd7,3'd7,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd4,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd5,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_30_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_29_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd5,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7},
'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd6,3'd6,3'd4,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6},
'{3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd6,3'd3,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd3,3'd2},
'{3'd6,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd1,3'd0},
'{3'd7,3'd6,3'd5,3'd4,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd6},
'{3'd3,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7},
'{3'd3,3'd3,3'd2,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd5},
'{3'd3,3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd2,3'd1,3'd0,3'd1,3'd2,3'd3,3'd6,3'd7,3'd7,3'd6,3'd5,3'd2,3'd1},
'{3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd2},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd6,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd4,3'd3,3'd3,3'd3,3'd4,3'd4,3'd5,3'd7},
'{3'd2,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd7},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd7},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd2,3'd3,3'd7},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd3,3'd7},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7},
'{3'd1,3'd2,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd5,3'd5,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7}};

parameter bit [2:0] SpriteTableR_29_30[31:0][31:0] = '{'{3'd5,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd3,3'd7,3'd6,3'd3,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7},
'{3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd3,3'd7},
'{3'd6,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd3,3'd7},
'{3'd4,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd3,3'd7},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd3,3'd7},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd5,3'd5,3'd4,3'd3,3'd2,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd4,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd7},
'{3'd1,3'd1,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7},
'{3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd7,3'd7,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd5,3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7},
'{3'd7,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd1,3'd5,3'd7},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd3,3'd1,3'd1,3'd2,3'd1,3'd5,3'd7},
'{3'd6,3'd6,3'd6,3'd5,3'd5,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd3,3'd0,3'd0,3'd1,3'd1,3'd5,3'd7},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd3,3'd0,3'd0,3'd1,3'd1,3'd6,3'd7},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd3,3'd0,3'd1,3'd1,3'd1,3'd6,3'd7},
'{3'd7,3'd7,3'd7,3'd4,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd1,3'd6,3'd7},
'{3'd7,3'd5,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd1,3'd6,3'd7},
'{3'd6,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd4,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd4,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7},
'{3'd3,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd4,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd4,3'd6,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd3,3'd1,3'd1,3'd0,3'd2,3'd7,3'd7},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd2,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd5,3'd5,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd6,3'd3,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd3,3'd5,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd3,3'd6,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd6,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd6,3'd6,3'd5,3'd3,3'd1,3'd2,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd6,3'd5,3'd7,3'd7}};

parameter bit [2:0] SpriteTableR_29_29[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd6,3'd3,3'd2,3'd6,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd6,3'd2,3'd1,3'd1,3'd5,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd6,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd2,3'd6,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd3,3'd6,3'd7,3'd6,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd3,3'd0,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd6},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd5,3'd3,3'd4,3'd7,3'd5,3'd2,3'd5,3'd7,3'd7,3'd7,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7},
'{3'd5,3'd4,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd1,3'd1,3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd6,3'd7},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd1,3'd0,3'd2,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd7},
'{3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd6,3'd5,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_29_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_28_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd5,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6,3'd5,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4},
'{3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd6,3'd6,3'd5,3'd5,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd2,3'd3,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd5,3'd6,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd1,3'd1,3'd3,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd1,3'd2,3'd3,3'd2,3'd2,3'd6,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd5,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd5,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd6,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd6,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd5,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_28_30[31:0][31:0] = '{'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd5,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0,3'd0},
'{3'd7,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd4,3'd5,3'd5,3'd4},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd2,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd7,3'd7,3'd4,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd7,3'd7,3'd4,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd4,3'd3,3'd2,3'd1,3'd2},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd6,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd4,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd6,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd7,3'd6,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd5,3'd2,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd5,3'd5,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd5,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd7,3'd7,3'd6,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd1,3'd1,3'd3,3'd7,3'd7,3'd7,3'd5,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd1,3'd1,3'd5,3'd7,3'd6,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd4,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd1,3'd3,3'd7,3'd5,3'd1,3'd1,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd1,3'd5,3'd7,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd4,3'd5},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd1,3'd6,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd6},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd2,3'd6,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd7,3'd6},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd3,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd5,3'd6,3'd6},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd3,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd6,3'd2,3'd6,3'd5},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd4,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd7,3'd7,3'd5,3'd7,3'd4},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd5,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd7,3'd6,3'd2},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd1,3'd5,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd7,3'd6,3'd3,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd2,3'd6,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd6,3'd4,3'd1,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd2,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd3,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd2,3'd1,3'd5,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_28_29[31:0][31:0] = '{'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd2,3'd2,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd6,3'd2,3'd3,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd1,3'd4,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd3,3'd1,3'd4,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd6},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd4,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd6,3'd7,3'd7},
'{3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd3,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd6,3'd6},
'{3'd2,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd1,3'd2,3'd7,3'd7,3'd4,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd3},
'{3'd4,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd2},
'{3'd7,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd5,3'd4,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd6,3'd6,3'd6,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_28_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_27_31[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7},
'{3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd5,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd4,3'd2,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd7},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd2,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd5,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd2,3'd5,3'd5,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd5,3'd5,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd6,3'd3,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd3,3'd1,3'd0,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd4,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd5,3'd1,3'd0,3'd1,3'd3,3'd1,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd6,3'd4,3'd0,3'd1,3'd4,3'd1,3'd0,3'd2,3'd6,3'd7,3'd7,3'd6,3'd3,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableR_27_30[31:0][31:0] = '{'{3'd1,3'd1,3'd0,3'd1,3'd2,3'd0,3'd0,3'd1,3'd4,3'd7,3'd3,3'd1,3'd5,3'd3,3'd2,3'd5,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd4,3'd6,3'd6,3'd6,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd4,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0},
'{3'd1,3'd2,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd5,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd5,3'd4,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd2,3'd3,3'd5,3'd6,3'd7},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd3,3'd4,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd6,3'd6,3'd5,3'd6,3'd5,3'd7,3'd5,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd6,3'd6,3'd3,3'd2,3'd5,3'd2,3'd5,3'd5,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd6,3'd3,3'd2,3'd5,3'd6,3'd2,3'd3,3'd5,3'd1,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd1,3'd1,3'd2,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd4,3'd2,3'd3,3'd6,3'd7,3'd6,3'd1,3'd1,3'd4,3'd2,3'd1,3'd5,3'd7,3'd7,3'd5,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd4,3'd7,3'd7,3'd4,3'd1,3'd0,3'd2,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd2,3'd3,3'd2,3'd5,3'd7,3'd7,3'd2,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd5,3'd7,3'd6,3'd2,3'd1,3'd1,3'd0,3'd1,3'd5,3'd7,3'd7,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd6,3'd1,3'd1,3'd0,3'd0,3'd2,3'd6,3'd7,3'd6,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd5,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd4,3'd6},
'{3'd2,3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd4,3'd6,3'd7,3'd7},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd3,3'd1,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd5,3'd7,3'd7,3'd7,3'd6},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0,3'd4,3'd7,3'd7,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd5,3'd3,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd1,3'd5,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd5,3'd5,3'd6},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd5,3'd1,3'd1,3'd0,3'd2,3'd6,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd5,3'd7,3'd7,3'd7,3'd6,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd4,3'd0,3'd1,3'd1,3'd5,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd4,3'd3,3'd2,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd4,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd6,3'd4,3'd1,3'd1,3'd3,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd1,3'd4,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_27_29[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd5,3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd6,3'd4,3'd1,3'd1,3'd4,3'd5,3'd6,3'd6,3'd5,3'd4,3'd4,3'd3,3'd4,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd4,3'd7,3'd6,3'd1,3'd0,3'd1,3'd1,3'd2,3'd3},
'{3'd7,3'd3,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd3,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7},
'{3'd7,3'd4,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd7,3'd5,3'd1,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd3,3'd5},
'{3'd6,3'd7,3'd5,3'd6,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd5,3'd7,3'd6,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd5,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd4,3'd2,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd3,3'd6},
'{3'd3,3'd7,3'd7,3'd6,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7},
'{3'd1,3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd7},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd6,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd3,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd6,3'd7,3'd7,3'd3,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd6,3'd7,3'd6,3'd3,3'd0,3'd0,3'd0,3'd3,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd6,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd6,3'd7,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_27_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd6,3'd7,3'd7,3'd7,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd1,3'd0,3'd2,3'd5,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd6,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd5,3'd3,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd7,3'd6,3'd7,3'd7,3'd7,3'd5,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd5,3'd7,3'd7,3'd7,3'd6,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd5,3'd7,3'd6,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd5,3'd5,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_26_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd6,3'd7,3'd7,3'd6,3'd4,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd4,3'd6,3'd4,3'd2,3'd4,3'd6,3'd4,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd7,3'd6,3'd4,3'd3,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd4,3'd6,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd3,3'd1,3'd2,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd5,3'd6,3'd6,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd3,3'd5,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd6,3'd6,3'd6,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd6,3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd0,3'd1,3'd2,3'd3,3'd5,3'd5,3'd6,3'd7,3'd7,3'd7,3'd5,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd5,3'd4,3'd2,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd6,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd7,3'd7,3'd5,3'd2,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd3,3'd3,3'd4,3'd6,3'd6,3'd5},
'{3'd0,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd2,3'd0,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd7},
'{3'd2,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd6,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd4,3'd6,3'd7,3'd4,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd2},
'{3'd2,3'd6,3'd6,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd6,3'd7,3'd7,3'd6,3'd4,3'd2},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd7,3'd7,3'd5},
'{3'd0,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7},
'{3'd0,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd1,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_26_30[31:0][31:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd5,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd5,3'd4,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd2,3'd1,3'd3,3'd7,3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd7,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd6,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd6,3'd7,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd7,3'd7},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd2,3'd2,3'd2,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd4,3'd7,3'd6,3'd1,3'd0,3'd1,3'd1,3'd2,3'd4,3'd5,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd6,3'd1,3'd2,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd5,3'd7,3'd5,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd5,3'd7,3'd5,3'd2,3'd4,3'd6,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6,3'd5,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7},
'{3'd3,3'd6,3'd5,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd4,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7},
'{3'd7,3'd7,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd3,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd7,3'd7,3'd7,3'd7},
'{3'd7,3'd7,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd2,3'd6,3'd7,3'd7,3'd6,3'd4},
'{3'd7,3'd7,3'd3,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd5,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0},
'{3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd0,3'd0},
'{3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd5,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd7,3'd7,3'd7,3'd6,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd5,3'd6,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd3,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd6,3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd7,3'd7,3'd5,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0,3'd1,3'd5,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd6,3'd7,3'd7,3'd7,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd1,3'd0,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_26_29[31:0][31:0] = '{'{3'd5,3'd7,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd4,3'd4,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd2,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd4,3'd3,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd4,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd6,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd7,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd2},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd7},
'{3'd7,3'd6,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd7,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7},
'{3'd7,3'd3,3'd4,3'd7,3'd7,3'd6,3'd4,3'd6,3'd7,3'd6,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd4,3'd2,3'd4,3'd5,3'd5,3'd5},
'{3'd3,3'd2,3'd6,3'd7,3'd7,3'd4,3'd1,3'd3,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd1,3'd2,3'd6,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd7,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd6,3'd7,3'd7,3'd4,3'd1,3'd1,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd7,3'd7,3'd6,3'd2,3'd1,3'd3,3'd5,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd4,3'd2,3'd5,3'd7,3'd7,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd6,3'd5,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd5,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd7,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_26_28[31:0][15:0] = '{'{3'd1,3'd1,3'd4,3'd7,3'd7,3'd7,3'd6,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd6,3'd4,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd3,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_25_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd6,3'd6,3'd5,3'd4,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd5,3'd7},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd5,3'd6,3'd7,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd5,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd1,3'd5},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd4,3'd5,3'd6,3'd6,3'd5,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd7},
'{3'd0,3'd1,3'd1,3'd2,3'd4,3'd6,3'd7,3'd5,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd5,3'd6,3'd7,3'd7,3'd7,3'd6,3'd2,3'd3,3'd4,3'd4,3'd4,3'd3,3'd1,3'd5,3'd7},
'{3'd1,3'd1,3'd3,3'd5,3'd7,3'd6,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd2,3'd3,3'd4,3'd3,3'd4,3'd2,3'd2,3'd7,3'd7},
'{3'd4,3'd5,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd2,3'd2,3'd4,3'd5,3'd7,3'd7,3'd7,3'd5,3'd4,3'd3,3'd4,3'd7,3'd4,3'd2,3'd3,3'd4,3'd4,3'd3,3'd2,3'd5,3'd7,3'd6},
'{3'd7,3'd5,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd5,3'd7,3'd7,3'd6,3'd5,3'd2,3'd1,3'd1,3'd1,3'd4,3'd6,3'd2,3'd2,3'd3,3'd4,3'd3,3'd1,3'd3,3'd7,3'd7,3'd3},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd6,3'd7,3'd7,3'd5,3'd3,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd5,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2,3'd6,3'd7,3'd5,3'd1},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd5,3'd6,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2,3'd6,3'd7,3'd5,3'd2,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd7,3'd4,3'd2,3'd3,3'd4,3'd3,3'd2,3'd5,3'd7,3'd6,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd6,3'd2,3'd3,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0},
'{3'd7,3'd6,3'd3,3'd2,3'd2,3'd2,3'd2,3'd4,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd6,3'd2,3'd3,3'd4,3'd3,3'd1,3'd4,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0,3'd0},
'{3'd6,3'd7,3'd7,3'd5,3'd2,3'd2,3'd2,3'd1,3'd3,3'd6,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd3,3'd6,3'd4,3'd2,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd7,3'd7,3'd6,3'd3,3'd2,3'd2,3'd1,3'd2,3'd6,3'd7,3'd5,3'd2,3'd1,3'd2,3'd6,3'd5,3'd2,3'd3,3'd3,3'd2,3'd2,3'd6,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd4,3'd2,3'd2,3'd2,3'd2,3'd5,3'd7,3'd5,3'd2,3'd5,3'd6,3'd2,3'd2,3'd4,3'd2,3'd2,3'd5,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd2,3'd4,3'd6,3'd7,3'd6,3'd3,3'd2,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd4,3'd2,3'd3,3'd3,3'd1,3'd4,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd7,3'd7,3'd4,3'd3,3'd2,3'd1,3'd3,3'd5,3'd4,3'd2,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd3,3'd6,3'd7,3'd6,3'd3,3'd1,3'd2,3'd1,3'd1,3'd3,3'd3,3'd2,3'd4,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_25_30[31:0][31:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd7,3'd4,3'd1,3'd2,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd3,3'd3,3'd2,3'd3,3'd6,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd7,3'd7,3'd3,3'd2,3'd3,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd5,3'd1,3'd3,3'd2,3'd2,3'd6,3'd7,3'd6,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd5,3'd2,3'd2,3'd2,3'd2,3'd6,3'd7,3'd6,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd5,3'd7,3'd6,3'd2,3'd2,3'd2,3'd2,3'd6,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd3,3'd3,3'd4,3'd6,3'd7,3'd7,3'd3,3'd1,3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd3,3'd1,3'd1,3'd0,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd3,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd6,3'd7,3'd7,3'd5,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd6,3'd7,3'd7,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd4,3'd2,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd3,3'd7,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd1,3'd5,3'd7,3'd7,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2,3'd3,3'd7,3'd7,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2,3'd2,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd6,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd6,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd5,3'd7,3'd7,3'd5,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd6,3'd7,3'd7,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd6,3'd6,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd1,3'd0,3'd1,3'd2,3'd3,3'd3,3'd4,3'd6,3'd7,3'd7},
'{3'd0,3'd0,3'd0,3'd1,3'd6,3'd7,3'd4,3'd4,3'd7,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd7,3'd7,3'd4,3'd2,3'd3,3'd4,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5},
'{3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd5,3'd6,3'd7,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd2},
'{3'd0,3'd0,3'd0,3'd2,3'd7,3'd7,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd5,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd7,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd4,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd6,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd6,3'd4,3'd2,3'd0,3'd1,3'd3,3'd7,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_25_29[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd6,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd6,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd0,3'd1,3'd5,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd5,3'd1,3'd0,3'd0,3'd1,3'd4,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd4,3'd6,3'd7,3'd7,3'd7,3'd6,3'd7,3'd7,3'd6,3'd1,3'd0,3'd1,3'd5,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd2,3'd5,3'd7,3'd7,3'd5,3'd4,3'd6,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd2,3'd1,3'd1,3'd3,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd7,3'd6,3'd5,3'd3,3'd2,3'd1,3'd0,3'd1,3'd0,3'd1,3'd4,3'd6,3'd7,3'd7,3'd7,3'd5,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd5,3'd5,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_25_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_24_31[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd2,3'd1,3'd0,3'd5,3'd2,3'd1,3'd7,3'd4,3'd1,3'd7,3'd5,3'd1,3'd7,3'd6,3'd1,3'd7,3'd4,3'd1,3'd6,3'd2,3'd1,3'd4,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_24_30[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd2,3'd1,3'd0,3'd4,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_24_29[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableR_24_28[2:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

logic [9:0] SpriteTableG;

parameter bit [7:0] SpritePaletteG[7:0] = '{8'd16, 8'd49, 8'd82, 8'd115, 8'd148, 8'd181, 8'd214, 8'd247};

	always_comb
	begin
		SpriteTableG = 10'd0;
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_31_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_31_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_31_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_31_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_30_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_30_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_30_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_30_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_29_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_29_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_29_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_29_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_28_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_28_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_28_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_28_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_27_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_27_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_27_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_27_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_26_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_26_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_26_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_26_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_25_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_25_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_25_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_25_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_24_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_24_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_24_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_24_28[Y_Index][X_Index];
		end
	end

parameter bit [2:0] SpriteTableG_31_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd3,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd4,3'd6,3'd6},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd4,3'd6,3'd6,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd5,3'd6,3'd6,3'd5,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd4,3'd6,3'd6,3'd5,3'd4,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_31_30[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd3,3'd5,3'd6,3'd6,3'd5,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd3,3'd5,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd5,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd5,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd4,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd4,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd3,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd2,3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd3,3'd1,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd2,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd2,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd2,3'd3,3'd3,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd2,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd2,3'd4,3'd1,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd3,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd1,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_31_29[31:0][31:0] = '{'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd2,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd4,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4,3'd2},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd4,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd4,3'd3,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd5,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd4,3'd4,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd4,3'd5,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd2},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd3,3'd2,3'd0,3'd1,3'd3,3'd3,3'd2,3'd3,3'd5,3'd6,3'd6},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd5,3'd6,3'd6,3'd5},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd4,3'd4,3'd3,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2},
'{3'd3,3'd4,3'd3,3'd2,3'd2,3'd4,3'd5,3'd6,3'd6,3'd6,3'd5,3'd5,3'd4,3'd3,3'd3,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd6,3'd6,3'd6,3'd5,3'd3,3'd1,3'd2},
'{3'd3,3'd3,3'd2,3'd4,3'd5,3'd6,3'd5,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd6,3'd5,3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0},
'{3'd6,3'd6,3'd5,3'd4,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd2,3'd3,3'd5,3'd6,3'd6,3'd5,3'd6,3'd6,3'd5,3'd3,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd6,3'd4,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd5,3'd4,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd5,3'd6,3'd6,3'd5,3'd3,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd6,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd4,3'd6,3'd3,3'd1,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_30_30[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd4,3'd3,3'd1,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd2,3'd0,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd3,3'd2,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd0,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd2,3'd4,3'd3,3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd4,3'd5,3'd4,3'd1,3'd2,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd5,3'd6,3'd6,3'd5,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd3,3'd2,3'd1,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd3,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd1,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd0,3'd0,3'd2,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd3,3'd3,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd3,3'd2,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd3,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd2,3'd0,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd3,3'd0,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_30_29[31:0][31:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd3,3'd4,3'd3,3'd3,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd4,3'd3,3'd1,3'd0,3'd2,3'd2,3'd1},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd1,3'd2},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd4,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd4,3'd3,3'd1,3'd2,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd3,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd4,3'd3,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd3,3'd3,3'd1},
'{3'd3,3'd1,3'd2,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd4,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd4,3'd2},
'{3'd0,3'd0,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd4,3'd5,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd3,3'd4},
'{3'd0,3'd1,3'd3,3'd1,3'd2,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2},
'{3'd0,3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd5,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd3,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd3,3'd1,3'd3,3'd4,3'd4,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd5,3'd4,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd5},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd5,3'd5,3'd5,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd5,3'd5,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd5,3'd5,3'd6,3'd6,3'd5,3'd5,3'd4,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd4,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd3,3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd5,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd3,3'd5,3'd5,3'd6,3'd6,3'd5,3'd4,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd2,3'd3,3'd5,3'd6,3'd6,3'd5,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2,3'd1,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0},
'{3'd3,3'd4,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd5,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd6,3'd5,3'd3,3'd2,3'd1,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd4,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd3,3'd5,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_29_30[31:0][31:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd3,3'd6,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd0,3'd0,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd3,3'd0,3'd1,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd2,3'd0,3'd1,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd2,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd0,3'd1,3'd0,3'd1,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd4},
'{3'd1,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd2,3'd3,3'd2,3'd3,3'd4,3'd3,3'd2,3'd1,3'd3,3'd4},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd2,3'd4,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd2,3'd2},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd2,3'd0,3'd1},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_29_29[31:0][31:0] = '{'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd4,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd4,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2},
'{3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd4,3'd4,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd4,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd4,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd0,3'd1,3'd2,3'd1,3'd1,3'd3,3'd4,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd5,3'd2,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd4,3'd5,3'd4,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd2,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd6,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4},
'{3'd2,3'd2,3'd3,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd6,3'd5,3'd6,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd1,3'd1},
'{3'd5,3'd5,3'd6,3'd6,3'd5,3'd5,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd5,3'd5,3'd4,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd5,3'd4,3'd1,3'd2,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd5,3'd5,3'd6,3'd5,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd4,3'd5,3'd6,3'd6,3'd6,3'd5,3'd5,3'd5,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd1,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd0,3'd1,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_28_30[31:0][31:0] = '{'{3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd1,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6},
'{3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd2,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd2,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd1,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd2,3'd4,3'd5,3'd6,3'd6,3'd5,3'd5,3'd5,3'd4,3'd2,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd1,3'd0,3'd1},
'{3'd2,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd2,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd1,3'd1},
'{3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd1,3'd1,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_28_29[31:0][31:0] = '{'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd3,3'd0,3'd1,3'd1,3'd0,3'd2,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd4,3'd2,3'd0,3'd1,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd5,3'd3,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd5,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd4,3'd4,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd3,3'd5,3'd4,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd3,3'd3,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd1,3'd2,3'd4,3'd5,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd4,3'd5,3'd4,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_31[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd5,3'd5,3'd5,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd4,3'd5,3'd5,3'd5,3'd4,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd4,3'd4,3'd5},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd2,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd5,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd4,3'd7,3'd5,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd5,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd5,3'd5,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd5,3'd5,3'd2,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd6,3'd2,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd3,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd4,3'd1,3'd1,3'd1,3'd3},
'{3'd2,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd6,3'd7,3'd5,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd5,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd7,3'd6,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd2,3'd6,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd5,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd6,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd5,3'd2,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1,3'd2,3'd5,3'd7,3'd7,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd4,3'd1,3'd1,3'd4,3'd2,3'd0,3'd2,3'd5,3'd7,3'd7,3'd7,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_27_30[31:0][31:0] = '{'{3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd4,3'd7,3'd3,3'd1,3'd5,3'd3,3'd2,3'd5,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd6,3'd6,3'd4,3'd6,3'd6,3'd5,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd4,3'd4,3'd5,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd6,3'd5,3'd5,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd7,3'd5,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd5,3'd7,3'd7,3'd7,3'd7,3'd7,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd5,3'd5,3'd5,3'd4,3'd1,3'd3,3'd6,3'd7,3'd5,3'd6,3'd5,3'd6,3'd5,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd6,3'd6,3'd3,3'd1,3'd4,3'd2,3'd5,3'd5,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd4,3'd6,3'd3,3'd1,3'd1,3'd3,3'd2,3'd2,3'd5,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6},
'{3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd1,3'd2,3'd1,3'd1,3'd3,3'd2,3'd1,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd6,3'd6,3'd6,3'd6,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd2,3'd1,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd3,3'd5,3'd3,3'd2,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6},
'{3'd6,3'd6,3'd6,3'd2,3'd1,3'd4,3'd5,3'd6,3'd3,3'd2,3'd2,3'd0,3'd0,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd4},
'{3'd6,3'd6,3'd5,3'd2,3'd4,3'd6,3'd6,3'd6,3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd4,3'd2,3'd1},
'{3'd6,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd6,3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd1,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd1,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd1,3'd0,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd0,3'd1,3'd2,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3,3'd1,3'd2,3'd3,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd4,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1,3'd2,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd4,3'd3,3'd3,3'd2,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd0,3'd0,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_27_29[31:0][31:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd2,3'd3,3'd1},
'{3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd2,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd4,3'd3},
'{3'd1,3'd2,3'd1,3'd2,3'd1,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd4,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd3,3'd1,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd3,3'd4,3'd3,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd3,3'd2,3'd1,3'd2,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1,3'd2,3'd2,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd4,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd3,3'd5,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd1,3'd2,3'd2,3'd3,3'd1,3'd1,3'd4,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_27_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd4,3'd2,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd2,3'd1,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd3,3'd5,3'd5,3'd5,3'd4,3'd3,3'd2,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd4,3'd5,3'd5,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd2,3'd1,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd4,3'd3,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd5,3'd4,3'd2,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd3,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd6,3'd7,3'd5,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd6,3'd6,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd4,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_26_30[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd6,3'd4,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd5,3'd6,3'd6,3'd4,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2},
'{3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd2,3'd3,3'd4,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2},
'{3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd6,3'd6,3'd6,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3},
'{3'd6,3'd5,3'd5,3'd3,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd2,3'd2,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd1,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd2,3'd1,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2},
'{3'd0,3'd1,3'd2,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd2,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd1,3'd2,3'd1,3'd3,3'd3,3'd4},
'{3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd4},
'{3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4},
'{3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_26_29[31:0][31:0] = '{'{3'd2,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd3,3'd3,3'd3,3'd4},
'{3'd1,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd4,3'd3,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd4,3'd2,3'd0,3'd1,3'd4,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd4,3'd4,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd2,3'd4,3'd4,3'd2,3'd2,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd2,3'd4,3'd5,3'd2,3'd1,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd5,3'd2,3'd0,3'd2,3'd3,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd4,3'd4,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd2,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd4,3'd3,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd1,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd2,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd1,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd2,3'd4,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd3,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd4,3'd2,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd2,3'd3,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd4,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd1,3'd4,3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd4,3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd3,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd4,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd4,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd4,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd3,3'd4,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd4,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd3,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd2,3'd4,3'd3,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_28[31:0][15:0] = '{'{3'd1,3'd1,3'd2,3'd4,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd5,3'd5,3'd5,3'd5,3'd5,3'd5,3'd4,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd5,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd4,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd2,3'd2,3'd3,3'd4,3'd6,3'd6,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd5,3'd6,3'd6,3'd6,3'd4,3'd2,3'd3,3'd1},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd4,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd6,3'd4,3'd2,3'd2,3'd2,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4,3'd6,3'd6,3'd5,3'd2,3'd2,3'd2,3'd0,3'd1},
'{3'd2,3'd2,3'd3,3'd5,3'd6,3'd6,3'd6,3'd5,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd5,3'd6,3'd5,3'd3,3'd2,3'd2,3'd1,3'd0,3'd1},
'{3'd4,3'd5,3'd5,3'd6,3'd6,3'd6,3'd4,3'd2,3'd2,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4,3'd6,3'd6,3'd4,3'd2,3'd2,3'd1,3'd0,3'd1,3'd0},
'{3'd4,3'd5,3'd6,3'd6,3'd6,3'd5,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd4,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd0},
'{3'd2,3'd3,3'd4,3'd5,3'd5,3'd2,3'd1,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4,3'd6,3'd5,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1,3'd2,3'd4,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd2,3'd3,3'd6,3'd5,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd4,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd5,3'd6,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd5,3'd6,3'd3,3'd1,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd4,3'd2,3'd1,3'd0,3'd2,3'd2,3'd3,3'd6,3'd4,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd5,3'd5,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd5,3'd5,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd5,3'd5,3'd2,3'd2,3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_30[31:0][31:0] = '{'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd4,3'd5,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd4,3'd5,3'd3,3'd2,3'd2,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd5,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd4,3'd3,3'd2,3'd3,3'd2,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd2,3'd4,3'd3,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd2,3'd1,3'd3,3'd3,3'd1,3'd2,3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd1,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd5,3'd5,3'd6,3'd6,3'd5,3'd4,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd2,3'd4,3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd1,3'd3,3'd3,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd4,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd2,3'd4,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd3,3'd3,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd3,3'd1,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd3,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd4,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd5,3'd3,3'd1,3'd0,3'd1,3'd0},
'{3'd4,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd5,3'd4,3'd4,3'd3,3'd2,3'd1,3'd2,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd4,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd4,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_29[31:0][31:0] = '{'{3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd2,3'd1,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd3,3'd3,3'd2,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd4,3'd4,3'd3,3'd4,3'd3,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd2,3'd4,3'd4,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_31[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd2,3'd0,3'd1,3'd2,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_30[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_29[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_28[2:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

logic [9:0] SpriteTableB;

parameter bit [7:0] SpritePaletteB[7:0] = '{8'd16, 8'd49, 8'd82, 8'd115, 8'd148, 8'd180, 8'd246, 8'd213};

	always_comb
	begin
		SpriteTableB = 10'd0;
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_31_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_31_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_31_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd992 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_31_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_30_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_30_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_30_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd960 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_30_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_29_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_29_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_29_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd928 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_29_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_28_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_28_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_28_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd896 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_28_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_27_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_27_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_27_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd864 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_27_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_26_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_26_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_26_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd832 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_26_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_25_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_25_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_25_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd800 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_25_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd992 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_24_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd960 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_24_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd928 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_24_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd768 && SpriteX < 10'd227 && SpriteY >= 10'd896 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_24_28[Y_Index][X_Index];
		end
	end

parameter bit [2:0] SpriteTableB_31_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_31_30[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableB_31_29[31:0][31:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_31_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_30_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableB_30_30[31:0][31:0] = '{'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd4,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_30_29[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_30_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_29_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd2,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0},
'{3'd2,3'd1,3'd1,3'd2,3'd4,3'd3,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2,3'd4,3'd5,3'd7,3'd4,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0}};

parameter bit [2:0] SpriteTableB_29_30[31:0][31:0] = '{'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd7,3'd6,3'd5,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd5,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4,3'd2,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd4,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd4,3'd3,3'd4,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_29_29[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_29_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_28_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableB_28_30[31:0][31:0] = '{'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableB_28_29[31:0][31:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_28_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_27_31[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd4,3'd5,3'd5,3'd4,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd6,3'd7,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd2,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd5,3'd5,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd3,3'd4,3'd2,3'd2,3'd5,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd5,3'd5,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd5,3'd5,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2,3'd5,3'd7,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd5,3'd7,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd7,3'd6,3'd3,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd2,3'd1,3'd2,3'd5,3'd6,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd5,3'd6,3'd5,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd7,3'd6,3'd5,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd1,3'd2,3'd2,3'd3,3'd2,3'd1,3'd2,3'd3,3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd7,3'd6,3'd7,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd4,3'd4,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2,3'd5,3'd6,3'd6,3'd3,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd5,3'd6,3'd6,3'd5,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd5,3'd6,3'd6,3'd7,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd5,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd5,3'd6,3'd6,3'd7,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd5,3'd5,3'd1,3'd1,3'd3,3'd2,3'd1,3'd2,3'd5,3'd6,3'd6,3'd7,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableB_27_30[31:0][31:0] = '{'{3'd4,3'd3,3'd3,3'd3,3'd4,3'd3,3'd2,3'd1,3'd3,3'd7,3'd3,3'd1,3'd4,3'd3,3'd2,3'd5,3'd6,3'd6,3'd6,3'd4,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd5,3'd7,3'd4,3'd7,3'd7,3'd5,3'd6,3'd6,3'd6,3'd4,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd3,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd7,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd7,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd2,3'd2,3'd3,3'd4,3'd4,3'd5,3'd7,3'd7,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd6,3'd5,3'd5,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd7,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd5,3'd6,3'd6,3'd6,3'd6,3'd6,3'd4,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd7,3'd7,3'd4,3'd5,3'd5,3'd7,3'd5,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd7,3'd7,3'd2,3'd1,3'd3,3'd2,3'd4,3'd5,3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd5,3'd2,3'd0,3'd0,3'd2,3'd2,3'd2,3'd5,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd3,3'd4,3'd2,3'd0,3'd1,3'd0,3'd1,3'd2,3'd1,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableB_27_29[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableB_27_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_26_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd5,3'd5,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd4,3'd3,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd0},
'{3'd5,3'd6,3'd6,3'd5,3'd4,3'd3,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd4,3'd7,3'd6,3'd4,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd4,3'd5,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableB_26_30[31:0][31:0] = '{'{3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd4,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableB_26_29[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_26_28[31:0][15:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_25_31[31:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_25_30[31:0][31:0] = '{'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_25_29[31:0][31:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_25_28[31:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_24_31[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_24_30[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_24_29[2:0][31:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableB_24_28[2:0][15:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

assign SpriteR = SpritePaletteR[SpriteTableR];
assign SpriteG = SpritePaletteG[SpriteTableG];
assign SpriteB = SpritePaletteB[SpriteTableB];

endmodule
